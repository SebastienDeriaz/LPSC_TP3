

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package colors_LUT is

    type colors_array is array (0 to 100) of std_logic_vector(7 downto 0);
    constant R : colors_array := ("00011100", "00011010", "00011000", "00010111", "00010110", "00010111", "00010111", "00011000", "00011010", "00011100", "00011110", "00100001", "00100100", "00101000", "00101100", "00110000", "00110101", "00111010", "00111111", "01000101", "01001010", "01010000", "01010110", "01011101", "01100011", "01101001", "01110000", "01110111", "01111110", "10000100", "10001011", "10010010", "10011001", "10100000", "10100110", "10101101", "10110011", "10111010", "11000000", "11000110", "11001100", "11010010", "11010111", "11011100", "11100001", "11100110", "11101010", "11101110", "11110010", "11110101", "11111000", "11111010", "11111100", "11111101", "11111110", "11111111", "11111110", "11111101", "11111100", "11111010", "11110111", "11110100", "11110000", "11101011", "11100101", "11011111", "11011000", "11010000", "11001000", "10111111", "10110110", "10101100", "10100010", "10011000", "10001110", "10000011", "01111001", "01101110", "01100100", "01011010", "01010000", "01000110", "00111100", "00110011", "00101011", "00100011", "00011100", "00010101", "00001111", "00001010", "00000110", "00000011", "00000001", "00000000", "00000000", "00000001", "00000011", "00000111", "00001101", "00010011", "00011100");
    constant G : colors_array := ("00100001", "00100100", "00101000", "00101100", "00110000", "00110100", "00111001", "00111110", "01000011", "01001000", "01001101", "01010011", "01011001", "01011110", "01100100", "01101010", "01110000", "01110110", "01111100", "10000011", "10001001", "10001111", "10010101", "10011011", "10100000", "10100110", "10101100", "10110001", "10110111", "10111100", "11000001", "11000101", "11001010", "11001110", "11010010", "11010110", "11011001", "11011100", "11011111", "11100001", "11100011", "11100100", "11100101", "11100110", "11100110", "11100110", "11100101", "11100100", "11100011", "11100001", "11011111", "11011101", "11011010", "11010111", "11010011", "11010000", "11001100", "11000111", "11000011", "10111110", "10111001", "10110011", "10101110", "10101000", "10100010", "10011100", "10010110", "10001111", "10001001", "10000010", "01111011", "01110100", "01101110", "01100111", "01100000", "01011001", "01010011", "01001101", "01000110", "01000000", "00111010", "00110101", "00101111", "00101010", "00100110", "00100001", "00011101", "00011010", "00010111", "00010100", "00010010", "00010000", "00001111", "00001110", "00001110", "00001111", "00010000", "00010010", "00010100", "00011000", "00011100");
    constant B : colors_array := ("01101011", "01101110", "01110010", "01110110", "01111010", "01111111", "10000011", "10001001", "10001110", "10010011", "10011001", "10011111", "10100101", "10101011", "10110000", "10110110", "10111100", "11000010", "11001000", "11001101", "11010011", "11011000", "11011101", "11100010", "11100110", "11101011", "11101110", "11110010", "11110101", "11111000", "11111010", "11111011", "11111101", "11111101", "11111101", "11111101", "11111100", "11111010", "11110111", "11110100", "11110000", "11101011", "11100101", "11011111", "11011000", "11010000", "11000111", "10111110", "10110100", "10101010", "10100000", "10010101", "10001011", "10000000", "01110101", "01101011", "01100000", "01010110", "01001100", "01000011", "00111010", "00110001", "00101001", "00100010", "00011100", "00010110", "00010010", "00001110", "00001011", "00001000", "00000110", "00000101", "00000100", "00000100", "00000100", "00000101", "00000110", "00001000", "00001001", "00001011", "00001101", "00010000", "00010010", "00010100", "00010111", "00011001", "00011100", "00011110", "00100000", "00100010", "00100100", "00100101", "00100110", "00100110", "00100111", "00100110", "00100101", "00100100", "00100010", "00011111", "00011100");

end package colors_LUT;
